module xorgate(x, y, z);
    input x, y;
    output z;

    assign z = x ^ y;
endmodule