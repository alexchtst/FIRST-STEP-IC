module hallo();

    initial begin
        $display("Hallo World");
        $finish;
    end

endmodule